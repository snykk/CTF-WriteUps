BZh91AY&SY�;�!  �߀Px���߰?���@��]��&��M�4�l�5=D�@��6�JhA"cQ��=F���M �L�j��=G��H�� h�#@ IiOҞI�<�b  ɓ@�*4ڃJI=�ťt?�Dh`���pmHM���:G�[�J��TI�zEn��h���m��S�RH����`J8d�-�e���{�$�'n��C�:�0ڼ�f�P�C�3�;fF�5��/5���PU5x�ey�%DgdgT�tjU��W�2�A=���; ��=h���/���l=�'��D�X�A�s�bS�����A��gk�!F���iG�y/��ٟ��;���㺃<������CK�^��,#F{f��GI�l^�xqpz"�V���Z��J�(�u�����+�bݤ��Eu�A���,�OC����Y����*�vfhߑ���ƞ����}o�@���dʙ^��7I@�����ȆJ���}x���:�,�M�d
6�;��#FKfL���֍S�Yr�kdϡcc�\R�mū�H̸��\�}7�K2y�Zn�|(9���3-<�0.��Lk��b�ё�L萊�E0���83�2
*�����f��r.��lf�ɋի��3�qX�h�+F<Ӏ�Z7m�����q:zj�v���Y3����[x���Yk��R��f��q9��]f�u9�i �(L���`u�֭�iӳ%]�wQ���=ml[9�w׳)��1S����z���a�Ơ�5)�+�6Z��1fG��Բ/�c�4H�Nf-�rE8P��;�!