BZh91AY&SYmW2 !߀Px���߰?���P���fU��%	�Sz��)�L�� � �h�&d`bba0�!�&�	&Bi�2z�J1��4i��&d`bba0�!�&�	"��'��I��dz� ���c@|`(p�� C�����bm����>��|�%V�s0�AVj_.�g�a��T�d}��d����H�	���|Lmo���<ֺ��EC���JFř�@����Mp~�PȊ.g�cvR���T�8-_���	B�W�\tR���d1w��k����h�u��D���y��2��ӹ��d�湎6?��܈�pC�S��.X�唱�MF:Fl�h���f5_��at$`֯*������n7ͨ{�~�DqG�eu���߲N>����!��[$E���y	�,��H�J��:qJ�|�)�(�=A��r�4�0�Z9�)��J���\�?~9F04�[+���K�C/�P�=l
��u�Wf%�U]<��F
��+�6�=�(����ǎ��Te�����4�,�g=��,'rƝH��l#h�$3�r*
��ds����ȵ^Y3��w����CJvc�RB�*��D�x�bD�p�4p���vz17f��9mm&*��Kj���)�Tر-�51*��ˠr���kc7끘2���
0Yʉ�#ۙ��Ad�a�$
Y�$�"]((�����k}��/P����A1[kP�ޠ�������Z�C��5nW�����i�. ��Č	��H�Xd��%�`���ł����i-�����s�ȻY�"e�lU�kJH����Cts4Z��Ө4�T8�=1�UA�x,/,w�a�fs��Į7	!��DE0��qN%�.�i�)Ϣ$��fJ����y@1��JV���"�(H6��� 